*Circuit Name
V1 VDD 0 2.5
M1 VDD N001 N001 VDD P_1u l=0.000046 w=0.000021
M2 VDD N001 N002 VDD P_1u l=0.000046 w=0.000021
M3 VDD N001 Vout VDD P_1u l=0.000046 w=0.000021
M4 N002 0 N004 N002 P_1u l=0.000008 w=0.000046
M5 N002 vi+ N003 N002 P_1u l=0.000008 w=0.000046
M6 N004 N004 VSS VSS N_1u l=0.000003 w=0.000015
M7 N003 N004 VSS VSS N_1u l=0.000003 w=0.000015
M8 Vout N003 VSS VSS N_1u l=0.000014 w=0.000025
C1 Vout N003 0.000000
I1 N001 VSS 0.000075
V2 VSS 0 -2.5
C2 0 Vout 1p
V3 Vi+ 0 AC 1
.model NMOS NMOS
.model PMOS PMOS
.ac oct 100 1 1meg
.include cmosedu_models.txt
.meas AC ganho FIND v(vout) AT 1
.end